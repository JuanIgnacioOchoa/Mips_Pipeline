library verilog;
use verilog.vl_types.all;
entity ALU is
    port(
        ALUOperation    : in     vl_logic_vector(3 downto 0);
        A               : in     vl_logic_vector(31 downto 0);
        B               : in     vl_logic_vector(31 downto 0);
        Shamt           : in     vl_logic_vector(4 downto 0);
        ProgramCounter  : in     vl_logic_vector(31 downto 0);
        bitLocForLoadAndSave: in     vl_logic_vector(15 downto 0);
        Zero            : out    vl_logic;
        NotZero         : out    vl_logic;
        JReg            : out    vl_logic;
        ALUResult       : out    vl_logic_vector(31 downto 0)
    );
end ALU;
